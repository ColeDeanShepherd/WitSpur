module mux4(
  input [3:0] in,
  input [1:0] select,
  output reg out
);
endmodule