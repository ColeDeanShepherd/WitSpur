module counter (
  input clock,
  input reset,
  output reg [3:0] out
);
  always @(posedge clock) begin
  end
endmodule