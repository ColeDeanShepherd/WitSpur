/*
Let's build a simple module which take two one-bit inputs, performs the "AND"
operation on the inputs, and outputs the resulting value.
*/

// First, let's declare an empty module named "my_AND".
module my_AND;
endmodule