/*
Let's build a half-adder: a simple module which takes two 1-bit input signals,
adds them, and outputs a "sum" bit (the least significant bit of the 2-bit sum)
and a "carry" bit (the most significant bit of the 2-bit sum).
*/

// First, let's declare an empty module named "half_adder".
module half_adder;
endmodule