module ram(
  input clock,
  input [7:0] address,
  output reg [7:0] data
);
endmodule